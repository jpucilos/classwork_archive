* Circuit netlist of NAND2 gate
* D Flip Flop Model
* jpucilos@stevens.edu 12/8/17
.include Mosis_tsmc_180nm.model

Vvdd VDD GND 3.3
VinA D GND dc 0 pulse 0 3.3 0ns 0.1ns 0.1ns 25ns 50ns
VinB CLK GND dc 0 pulse 0 3.3 12ns 0.1ns 0.1ns 25ns 50ns


*Invert D - output inv
Invert1 inv D GND GND NMOS L=0.18um W=0.8um
Invert2 inv D VDD VDD PMOS L=0.18um W=0.8um

*NAND Gate for D and Clk - output W
MN11 A1 D GND GND NMOS L=0.18um W=0.8um
MN12 W CLK A1 GND NMOS L=0.18um W=0.8um
MP11 W D VDD VDD PMOS L=0.18um W=0.8um
MP12 W CLK VDD VDD PMOS L=0.18um W=0.8um
Cout1 W GND 100fF

*NAND Gate for inv and Clk - output X
MN21 A2 inv GND GND NMOS L=0.18um W=0.8um
MN22 X CLK A2 GND NMOS L=0.18um W=0.8um
MP21 X inv VDD VDD PMOS L=0.18um W=0.8um
MP22 X CLK VDD VDD PMOS L=0.18um W=0.8um
Cout2 X GND 100fF

*NAND Gate for W and Y - output Q
MN31 A3 W GND GND NMOS L=0.18um W=0.8um
MN32 Q Y A3 GND NMOS L=0.18um W=0.8um
MP31 Q W VDD VDD PMOS L=0.18um W=0.8um
MP32 Q Y VDD VDD PMOS L=0.18um W=0.8um
Cout3 Q GND 100fF

*NAND Gate for X and Z - output Y
MN41 A4 X GND GND NMOS L=0.18um W=0.8um
MN42 Y Q A4 GND NMOS L=0.18um W=0.8um
MP41 Y X VDD VDD PMOS L=0.18um W=0.8um
MP42 Y Q VDD VDD PMOS L=0.18um W=0.8um
Cout4 Y GND 100fF

.tran .1ns 100ns



* D Flip Flop Model - Master Slave Configuration
* jpucilos@stevens.edu 12/8/17
.include Mosis_tsmc_180nm.model
*
Vvdd VDD GND 3.3
VinD D GND dc 0 pulse 0 3.3 0ns 0.1ns 0.1ns 25ns 50ns
VinInv inv GND dc 0 pulse 0 3.3 25ns 0.1ns 0.1ns 25ns 50ns
VinClk CLK GND dc 0 pulse 0 3.3 12ns 0.1ns 0.1ns 25ns 50ns
*
.subckt NAND A B C
M1 S A GND GND NMOS L=0.18um W=0.8um
M2 C B S GND NMOS L=0.18um W=0.8um
M3 C A VDD VDD PMOS L=0.18um W=0.8um
M4 C B VDD VDD PMOS L=0.18um W=0.8um
Cout C GND 100fF
.ends
*
* Master
*
X1 D CLK W NAND
X2 inv CLK X NAND
X3 W Q_bar Q NAND
X4 X Q Q_bar NAND
*
.tran .1ns 100ns



* Circuit netlist of NAND2 gate
* D Flip Flop Model
* jpucilos@stevens.edu 12/8/17
.include Mosis_tsmc_180nm.model

Vvdd VDD GND 3.3
VinA D GND dc 0 pulse 0 3.3 0ns 0.1ns 0.1ns 25ns 50ns
VinB CLK GND dc 0 pulse 0 3.3 12ns 0.1ns 0.1ns 25ns 50ns
VinInv inv GND dc 0 pulse 0 3.3 25ns 0.1ns 0.1ns 25ns 50ns

*NAND Gate for D and Clk - output W
MN11 A1 D GND GND NMOS L=0.18um W=0.8um
MN12 W CLK A1 GND NMOS L=0.18um W=0.8um
MP11 W D VDD VDD PMOS L=0.18um W=0.8um
MP12 W CLK VDD VDD PMOS L=0.18um W=0.8um
Cout1 W GND 100fF

*NAND Gate for inv and Clk - output X
MN21 A2 inv GND GND NMOS L=0.18um W=0.8um
MN22 X CLK A2 GND NMOS L=0.18um W=0.8um
MP21 X inv VDD VDD PMOS L=0.18um W=0.8um
MP22 X CLK VDD VDD PMOS L=0.18um W=0.8um
Cout2 X GND 100fF

*NAND Gate for W and Y - output Q
MN31 A3 W GND GND NMOS L=0.18um W=0.8um
MN32 Q Y A3 GND NMOS L=0.18um W=0.8um
MP31 Q W VDD VDD PMOS L=0.18um W=0.8um
MP32 Q Y VDD VDD PMOS L=0.18um W=0.8um
Cout3 Q GND 100fF

*NAND Gate for X and Z - output Y
MN41 A4 X GND GND NMOS L=0.18um W=0.8um
MN42 Y Q A4 GND NMOS L=0.18um W=0.8um
MP41 Y X VDD VDD PMOS L=0.18um W=0.8um
MP42 Y Q VDD VDD PMOS L=0.18um W=0.8um
Cout4 Y GND 100fF

.tran .1ns 100ns



* D Flip Flop Model - Master Slave Configuration
* jpucilos@stevens.edu 12/8/17
.include Mosis_tsmc_180nm.model
*
Vvdd VDD GND 3.3
VinD D GND dc 0 pulse 0 3.3 0ns 0.1ns 0.1ns 25ns 50ns
VinClk CLK GND dc 0 pulse 0 3.3 12ns 0.1ns 0.1ns 25ns 50ns
*
.subckt NAND A B Y
MN1 X A GND GND NMOS L=0.18um W=0.8um
MN2 Y B X GND NMOS L=0.18um W=0.8um
MP1 Y A VDD VDD PMOS L=0.18um W=0.8um
MP2 Y B VDD VDD PMOS L=0.18um W=0.8um
Cout Y GND 100fF
.ends
*
* Master
*
* Invert D - output inv
MInv1 inv D GND GND NMOS L=0.18um W=0.8um
MInv2 inv D VDD VDD PMOS L=0.18um W=0.8um
*

X1 W CLK D NAND
*X2 inv CLK X NAND
*X3 W Q_bar Q NAND
*X4 X Q Q_bar NAND
*
.tran .1ns 100ns
.end



